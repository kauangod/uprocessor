library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity rom is
  port (
    clk     : in std_logic;
    address : in unsigned(6 downto 0)   := (others => '0');
    data    : out unsigned(16 downto 0) := (others => '0')
  );
end entity;

architecture a_rom of rom is
    type mem is array (0 to 127) of unsigned(16 downto 0);
    constant rom_content : mem := (
      0  => B"0000000000_111_0001", --LD A,0
      1  => B"0000000000_000_0001", --LD R0,0
      2  => B"0000000001_001_0001", --LD R1,1
      3  => B"0000000101_010_0001", --LD R2,5

      4  => B"0000_000_100_111_0010", --MOV A,R0
      5  => B"0000_001_000_111_0010", --ADD R1
      6  => B"0000_111_100_000_0010", --MOV R0,A
      7  => B"0000_111_111_000_0010", --SW A,R0
      8  => B"0000_010_011_111_0010", --SRLI R2
      9  => B"0000000_001_000_0011", --CMPI 0
      10 => B"1111010_010_000_0011", --BLE -6

      11 => B"0000000010_000_0001", --LD 2,R0
      12 => B"0000000010_001_0001", --LD 2,R1

      13 => B"0000_000_100_111_0010", --MOV A,R0
      14 => B"0000_001_000_111_0010", --ADD R1 
      15 => B"0000_111_100_000_0010", --MOV R0,A
      16 => B"0000000000_111_0001", --LD A,0
      17 => B"0000_111_111_000_0010", --SW A,R0
      18 => B"0000_000_100_111_0010", --MOV A,R0
      19 => B"0000_010_011_111_0010", --SRLI R2
      20 => B"0000000_001_000_0011", --CMPI 0
      21 => B"1111000_010_000_0011", --BLE -8

      22 => B"0000000011_000_0001", --LD 3,R0
      23 => B"0000000011_001_0001", --LD 3,R1

      24 => B"0000_000_100_111_0010", --MOV A,R0
      25 => B"0000_001_000_111_0010", --ADD R1
      26 => B"0000_111_100_000_0010", --MOV R0,A
      27 => B"0000000000_111_0001", --LD A,0
      28 => B"0000_111_111_000_0010", --SW A,R0
      29 => B"0000_000_100_111_0010", --MOV A,R0
      30 => B"0000_010_011_111_0010", --SRLI R2
      31 => B"0000000_001_000_0011", --CMPI 0
      32 => B"1111000_010_000_0011", --BLE -8

      33 => B"0000000101_000_0001", --LD 5,R0
      34 => B"0000000101_001_0001", --LD 5,R1

      35 => B"0000_000_100_111_0010", --MOV A,R0
      36 => B"0000_001_000_111_0010", --ADD R1
      37 => B"0000_111_100_000_0010", --MOV R0,A
      38 => B"0000000000_111_0001", --LD A,0
      39 => B"0000_111_111_000_0010", --SW A,R0
      40 => B"0000_000_100_111_0010", --MOV A,R0
      41 => B"0000_010_011_111_0010", --SRLI R2
      42 => B"0000000_001_000_0011", --CMPI 0
      43 => B"1111000_010_000_0011", --BLE -8

      44 => B"0000000001_000_0001", --LD 1,R0
      45 => B"0000000001_001_0001", --LD 1,R1

      46 => B"0000_000_100_111_0010", --MOV A,R0
      47 => B"0000_001_000_111_0010", --ADD R1
      48 => B"0000_111_100_000_0010", --MOV R0,A
      49 => B"0000_000_110_111_0010", --LW A,R0
      50 => B"0000_111_100_110_0010", --MOV R6,A
      51 => B"0000_000_100_111_0010", --MOV A,R0
      52 => B"0000_010_011_111_0010", --SRLI R2
      53 => B"0000000_001_000_0011", --CMPI 0
      54 => B"1111000_010_000_0011", --BLE -8

      others => (others => '0')
    );

begin
    process (clk)
    begin
      if (rising_edge(clk)) then
        data <= rom_content(to_integer(address));
      end if;
    end process;
end architecture;