library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity rom is
  port (
    clk     : in std_logic;
    address : in unsigned(6 downto 0)   := (others => '0');
    data    : out unsigned(16 downto 0) := (others => '0')
  );
end entity;

architecture a_rom of rom is
    type mem is array (0 to 127) of unsigned(16 downto 0);
    constant rom_content : mem := (
      0  => B"0000000000_111_0001", --ld 0 A
      1  => B"0000000000_000_0001", --ld 0 r0
      2  => B"0000000001_001_0001", --ld 1 r1
      3  => B"0000000101_010_0001", --ld 5 r2

      4  => B"0000_000_100_111_0010", --mov r0 A   
      5  => B"0000_001_000_111_0010", --add A, r1
      6  => B"0000_111_100_000_0010", --mov A r0            
      7  => B"0000_111_111_000_0010", --sw A, r0 - insert
      8  => B"0000_010_011_111_0010", --slr r2
      9  => B"0000000_001_000_0011", --cmpi 0 
      10 => B"1111010_010_000_0011", --ble -6 (insert)

      11 => B"0000000010_000_0001", --ld 2 r0
      12 => B"0000000010_001_0001", --ld 2 r1

      13 => B"0000_000_100_111_0010", --mov r0 A - loop2   
      14 => B"0000_001_000_111_0010", --add A, r1
      15 => B"0000_111_100_000_0010", --mov A r0  
      16 => B"0000000000_111_0001", --ld 0 A          
      17 => B"0000_111_111_000_0010", --sw A, r0
      18 => B"0000_000_100_111_0010", --mov r0 A
      19 => B"0000_010_011_111_0010", --slr r2
      20 => B"0000000_001_000_0011", --cmpi 0 
      21 => B"1111000_010_000_0011", --ble -8 (loop2)

      22 => B"0000000011_000_0001", --ld 3 r0
      23 => B"0000000011_001_0001", --ld 3 r1

      24 => B"0000_000_100_111_0010", --mov r0 A - loop2   
      25 => B"0000_001_000_111_0010", --add A, r1
      26 => B"0000_111_100_000_0010", --mov A r0  
      27 => B"0000000000_111_0001", --ld 0 A          
      28 => B"0000_111_111_000_0010", --sw A, r0
      29 => B"0000_000_100_111_0010", --mov r0 A
      30 => B"0000_010_011_111_0010", --slr r2
      31 => B"0000000_001_000_0011", --cmpi 0 
      32 => B"1111000_010_000_0011", --ble -8 (loop2)

      33 => B"0000000101_000_0001", --ld 5 r0
      34 => B"0000000101_001_0001", --ld 5 r1

      35 => B"0000_000_100_111_0010", --mov r0 A - loop2   
      36 => B"0000_001_000_111_0010", --add A, r1
      37 => B"0000_111_100_000_0010", --mov A r0  
      38 => B"0000000000_111_0001", --ld 0 A          
      39 => B"0000_111_111_000_0010", --sw A, r0
      40 => B"0000_000_100_111_0010", --mov r0 A
      41 => B"0000_010_011_111_0010", --slr r2
      42 => B"0000000_001_000_0011", --cmpi 0 
      43 => B"1111000_010_000_0011", --ble -8 (loop2)

      44 => B"0000000000_000_0001", --ld 0 r0
      45 => B"0000000001_001_0001", --ld 1 r1

      46 => B"0000_000_100_111_0010", --mov r0 A - leitura
      47 => B"0000_001_000_111_0010", --add A r1
      48 => B"0000_111_100_000_0010", --mov A r0
      49 => B"0000_000_110_111_0010", --lw A r0
      50 => B"0000_111_100_110_0010", --mov A r6
      51 => B"0000_000_100_111_0010", --mov r0 A
      52 => B"0000_010_011_111_0010", --slr r2
      53 => B"0000000_001_000_0011", --cmpi 0 
      54 => B"1111000_010_000_0011", --ble -8 (insert)

      others => (others => '0')
    );

begin
    process (clk)
    begin
      if (rising_edge(clk)) then
        data <= rom_content(to_integer(address));
      end if;
    end process;
end architecture;